`timescale 1ns/1ps

module tb_asynch_fifo;
    logic clk_w;
    logic rst_w;